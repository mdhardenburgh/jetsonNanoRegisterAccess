module mainTop();

endmodule
